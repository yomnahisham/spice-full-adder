
.include ./MOSFET_models_0p5_0p18-3.inc
.include ./subcircuits.cir


VDD p_s 0 DC 1.8


VA A 0 PULSE(0 1.8 1n 1p 1p 40n 80n)
VB B 0 PULSE(0 1.8 2n 1p 1p 20n 40n)
VCi Ci 0 PULSE(0 1.8 4n 1p 1p 10n 20n)


* G1: XNOR(A,B)
XX1 p_s A B x1 0 XNOR Wn=0.143u Wp=0.286u
* G2: INV
XI1 p_s x1 x1_inv 0 INVERTER Wn=0.226u Wp=0.452u
* G3: XNOR(x1_inv, Ci)
XX2 p_s x1_inv Ci x2 0 XNOR Wn=0.357u Wp=0.714u
* G4: INV
XI2 p_s x2 x2_inv 0 INVERTER Wn=0.567u Wp=1.134u
* G5: OUT buffer INV
XI3 p_s x2_inv S_buf 0 INVERTER Wn=0.9u Wp=1.8u
* G6: Final output INV (corrects inversion from buffer)
XI4 p_s S_buf S 0 INVERTER Wn=0.9u Wp=1.8u

XNA1 p_s A B nab 0 NAND Wn=0.226u Wp=0.452u
XIA1 p_s nab ab 0 INVERTER Wn=0.357u Wp=0.714u

XNA2 p_s x1_inv Ci ncix 0 NAND Wn=0.226u Wp=0.452u
XIA2 p_s ncix cix 0 INVERTER Wn=0.357u Wp=0.714u

XNO p_s ab cix nor_out 0 NOR Wn=0.567u Wp=1.134u
XIO p_s nor_out Co 0 INVERTER Wn=0.9u Wp=1.8u

RloadS S S_load 1k
CloadS S_load 0 0.2p
RloadCo Co Co_load 1k
CloadCo Co_load 0 0.2p


.meas tran tPLH_S TRIG V(A) VAL=0.9 RISE=1 TARG V(S) VAL=0.9 RISE=1
.meas tran tPHL_S TRIG V(Ci) VAL=0.9 FALL=1 TARG V(S) VAL=0.9 FALL=1 TD=13n
.meas tran tPLH_C TRIG V(B) VAL=0.9 RISE=1 TARG V(Co) VAL=0.9 RISE=1
.meas tran tPHL_C TRIG V(B) VAL=0.9 FALL=1 TARG V(Co) VAL=0.9 FALL=1


.meas tran Etotal INTEG -V(p_s)*I(VDD) FROM=0 TO=80n
.meas tran Pavg PARAM='Etotal/80n'

.tran 85n

.plot v(S) v(Co) v(A) v(B) v(Ci) -I(VDD)

.end
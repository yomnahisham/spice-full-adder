* 		Level-1 Model for PMOS in model 0.18um CMOS Technology
.model PMOS0P18	PMOS(Level=1 VTO=-0.5 GAMMA=0.3 PHI=0.8
+		LD=10E-09 WD=0 UO=100 LAMBDA=0.17 TOX=4.08E-9 PB=0.9 CJ=1E-3
+		CJSW=2.04E-10 MJ=0.45 MJSW=0.29 CGDO=3.43E-10 JS=4.0E-7 CGBO=3.5E-10
+		CGSO=3.43E-10)


* 		Level-1 Model for NMOS in model 0.18um CMOS Technology
.model NMOS0P18	NMOS(Level=1 VTO=0.5 GAMMA=0.3 PHI=0.84
+		LD=10E-09 WD=0 UO=450 LAMBDA=0.2 TOX=4.08E-9 PB=0.9 CJ=1.6E-3
+		CJSW=2.04E-10 MJ=0.5 MJSW=0.2 CGDO=3.67E-10 JS=8.38E-6 CGBO=3.8E-10
+		CGSO=3.67E-10)

.subckt INVERTER VDD A Y Ground
MP Y A VDD VDD PMOS0P18 w=1.8u l=0.18u
MN Y A Ground Ground NMOS0P18 w=0.9u l=0.18u
.ends INVERTER



.subckt XNOR VDD A B Y Ground

XInverter1 VDD A A_n 0 INVERTER
XInverter2 VDD B B_n 0 INVERTER

MP1 wire_1 B_n VDD VDD PMOS0P18 w=1.8u l=0.18u
MP2 wire_1 A VDD VDD PMOS0P18 w=1.8u l=0.18u

MP3 Y B wire_1 wire_1 PMOS0P18 w=1.8u l=0.18u
MP4 Y A_n wire_1 wire_1 PMOS0P18 w=1.8u l=0.18u

MN1 Y B_n wire_2 wire_2 NMOS0P18 w=0.9u l=0.18u
MN2 wire_2 A Ground Ground NMOS0P18 w=0.9u l=0.18u

MN3 Y B wire_3 wire_3 NMOS0P18 w=0.9u l=0.18u
MN4 wire_3 A_n Ground Ground NMOS0P18 w=0.9u l=0.18u
.ends XNOR



.subckt NOR VDD A B Y Ground
MP1 wire_1 A VDD VDD PMOS0P18 w=1.8u l=0.18u
MP2 Y B wire_1 wire_1 NMOS0P18 w=1.8u l=0.18u

MN1 Y A Ground Ground NMOS0P18 w=0.9u l=0.18u
MN2 Y B Ground Ground NMOS0P18 w=0.9u l=0.18u
.ends NOR



.subckt NAND VDD A B Y Ground
MP1 Y B VDD VDD PMOS0P18 w=1.8u l=0.18u
MP2 Y A VDD VDD PMOS0P18 w=1.8u l=0.18u

MN1 Y B wire wire NMOS0P18 w=0.9u l=0.18u
MN2 wire A Ground Ground NMOS0P18 w=0.9u l=0.18u
.ends NAND

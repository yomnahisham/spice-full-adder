
.include ./MOSFET_models_0p5_0p18-3.inc
.include ./subcircuits.cir

* Full adder truth table via DC operating point; step A,B,Ci over {0,1}
VDD vdd 0 DC 1.8

* DC inputs (driven by stepped params)
.param A=0 B=0 Ci=0
VA A 0 DC {A}
VB B 0 DC {B}
VCi Ci 0 DC {Ci}

* Instantiate same gates and sizing as in full_adder_opt.cir
XX1 vdd A B xnor1 0 XNOR Wn=0.143u Wp=0.286u
XI1 vdd xnor1 xor1 0 INVERTER Wn=0.226u Wp=0.452u
XX2 vdd xor1 Ci xnor2 0 XNOR Wn=0.357u Wp=0.714u
XI2 vdd xnor2 S 0 INVERTER Wn=0.567u Wp=1.134u

XNA1 vdd A B nab 0 NAND Wn=0.226u Wp=0.452u
XIA1 vdd nab ab 0 INVERTER Wn=0.357u Wp=0.714u
XNA2 vdd xor1 Ci nci_xor1 0 NAND Wn=0.226u Wp=0.452u
XIA2 vdd nci_xor1 ci_xor1 0 INVERTER Wn=0.357u Wp=0.714u
XNO vdd ab ci_xor1 nor_out 0 NOR Wn=0.567u Wp=1.134u
XIO vdd nor_out Co 0 INVERTER Wn=0.9u Wp=1.8u

* Loads to match full_adder_opt.cir
RloadS S S_load 1k
CloadS S_load 0 0.2p
RloadCo Co Co_load 1k
CloadCo Co_load 0 0.2p

* Step the inputs through all combinations
.step param A list 0 1
.step param B list 0 1
.step param Ci list 0 1

* Operating point and print outputs (one line per step)
.op
.print dc V(A) V(B) V(Ci) V(S) V(Co)

.end


.include ./MOSFET_models_0p5_0p18-3.inc
VDD p_s 0 DC 3.3
Vin g 0 DC 1m
.DC Vin 0 3.3 1m

Rld m load 1k

Cld load 0 0.5p

* Matched design: PMOS W = NMOS W = 1.25u
MP m g p_s p_s PMOS0P5 w=1.25u l=0.5u
MN m g 0 0 NMOS0P5 w=1.25u l=0.5u

.end